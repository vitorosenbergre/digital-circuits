library verilog;
use verilog.vl_types.all;
entity BinDec_vlg_vec_tst is
end BinDec_vlg_vec_tst;
