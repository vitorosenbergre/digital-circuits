library verilog;
use verilog.vl_types.all;
entity demux8x1_vlg_vec_tst is
end demux8x1_vlg_vec_tst;
