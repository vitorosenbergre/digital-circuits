library verilog;
use verilog.vl_types.all;
entity cicuitoAtividade1_vlg_vec_tst is
end cicuitoAtividade1_vlg_vec_tst;
